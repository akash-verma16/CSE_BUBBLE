//! CS220 Assignment 7
//! Devansh Kumar Jha 200318
//! Shivang Pandey 200941

//! These are the memory modules which will be called and used in the processor module. They all will be present in the
//! write mode until the loading phase of the processor is running after that instruction memory would convert into
//! read only mode but the data memory would still be present in write mode to the user.

/// This is the module which will be used as the source of memory and this has the following controls as explained
// clk - The synchronizing signal for all the phases of the processor machine.
// reset - The reset signal to delete and restart the whole memory.
// in - The data which is send as input for storing in memory.
// out - The data which is being asked for from memory.
// mode - The working mode of the memory currently. 0 means write mode and 1 means read only mode.
// address_a - The address at which the input is filled by the memory.
// address_b - The address from which output is generated by the memory.
// writeEnable - In write mode when we have to refrain from writing into memory disable this flag.
module veda_instruction #(parameter width = 32, parameter depth = 256, parameter len = 8, parameter start = 0) (
    clk,reset,
    in,out,mode,address_a,address_b,
    writeEnable
);
    input wire [width-1:0] in;
    input wire [len-1:0] address_a,address_b;
    input wire clk,reset,mode,writeEnable;                                // Mode 0 means write mode and Mode 1 means read mode
    output wire [width-1:0] out;
    
    reg [width-1:0] memory[0:depth-1];
    reg [width-1:0] dataout,cur;
    integer i;

    // Setting the memory at erased state.
    initial begin
        if(start == 0) begin cur <= 0; end
    end

    // Load the default program of bubble sort if start is set to HIGH.
    initial begin
        if(start == 1) begin
            // Write program to enter instruction memory into the machine
            memory[0]  <= 32'b001000_00110_11011_0000000000001010;               // lw $27, 10($6)  $s3 = 10 (main)
            memory[1]  <= 32'b000001_00110_11010_0000000000001011;               // addi $26, $6, 11  $s2 = 11
            memory[2]  <= 32'b000001_00110_01001_0000000000000010;               // addi $9, $6, 2
            memory[3]  <= 32'b010010_00000000000000000000100000;                 // jal 32
            memory[4]  <= 32'b010010_00000000000000000000001001;                 // jal 9
            memory[5]  <= 32'b000001_00110_01001_0000000000000110;               // addi $9, $6, 6
            memory[6]  <= 32'b010010_00000000000000000000100000;                 // jal 32
            memory[7]  <= 32'b000001_00110_01000_0000000000000010;               // addi $8, $6, 2
            memory[8]  <= 32'b010101_00000000000000000000000000;                 // syscall
            memory[9]  <= 32'b000001_00110_10001_0000000000000000;               // addi $17, $6, 0 (bubble_sort)
            memory[10] <= 32'b000000_11011_10001_10010_00000_000001;             // sub $18, $27, $17 (outer)
            memory[11] <= 32'b000001_10010_10010_1111111111111111;               // addi $18, $18, -1
            memory[12] <= 32'b000001_00110_10011_0000000000000000;               // addi $19, $6, 0
            memory[13] <= 32'b000000_10011_10010_11001_00000_000001;             // sub $25, $19, $18
            memory[14] <= 32'b010011_11001_00110_11111_00000_000000;             // slt $31, $25, $6
            memory[15] <= 32'b001010_00110_11111_0000000000001101;               // beq $31, $6, 13
            memory[16] <= 32'b001101_00110_11001_0000000000001100;               // bgte $25, $6, 12
            memory[17] <= 32'b000111_00000_10011_10100_00000_000000;             // sll $20, $19, 0 (inner)
            memory[18] <= 32'b000000_10100_11010_10100_00000_000000;             // add $20, $20, $26
            memory[19] <= 32'b000001_10100_10101_0000000000000001;               // addi $21, $20, 1
            memory[20] <= 32'b001000_10100_10110_0000000000000000;               // lw $22, 0($20)
            memory[21] <= 32'b001000_10101_10111_0000000000000000;               // lw $23, 0($21)
            memory[22] <= 32'b000000_10110_10111_11000_00000_000001;             // sub $24, $22, $23
            memory[23] <= 32'b010011_11000_00110_11111_00000_000000;             // slt $31, $24, $6
            memory[24] <= 32'b001011_00110_11111_0000000000000010;               // bne $31, $6, 2
            memory[25] <= 32'b001001_10101_10110_0000000000000000;               // sw $22, 0($21)
            memory[26] <= 32'b001001_10100_10111_0000000000000000;               // sw $23, 0($20)
            memory[27] <= 32'b000001_10011_10011_0000000000000001;               // addi $19, $19, 1 (inend)
            memory[28] <= 32'b001011_10010_10011_1111111111110100;               // bne $19, $18, -12
            memory[29] <= 32'b000001_10001_10001_0000000000000001;               // addi $17, $17, 1 (oend)
            memory[30] <= 32'b001011_11011_10001_1111111111101011;               // bne $17, $27, -21
            memory[31] <= 32'b010001_00000000000000000000010000;                 // jr $16 (end1)
            memory[32] <= 32'b000001_00110_01000_0000000000000111;               // addi $8, $6, 7 (print)
            memory[33] <= 32'b000001_01001_01010_0000000000000000;               // addi $10, $9, 0
            memory[34] <= 32'b001000_01010_01010_0000000000000000;               // lw $10, 0($10)
            memory[35] <= 32'b000001_01001_01011_0000000000000001;               // addi $11, $9, 1
            memory[36] <= 32'b001000_01011_01011_0000000000000000;               // lw $11, 0($11)
            memory[37] <= 32'b000001_01001_01100_0000000000000010;               // addi $12, $9, 2
            memory[38] <= 32'b001000_01100_01100_0000000000000000;               // lw $12, 0($12)
            memory[39] <= 32'b000001_01001_01101_0000000000000011;               // addi $13, $9, 3
            memory[40] <= 32'b001000_01101_01101_0000000000000000;               // lw $13, 0($13)
            memory[41] <= 32'b010101_00000000000000000000000000;                 // syscall
            memory[42] <= 32'b000001_00110_10010_0000000000000000;               // addi $18, $6, 0
            memory[43] <= 32'b000001_11010_10001_0000000000000000;               // addi $17, $26, 0
            memory[44] <= 32'b000001_00110_01000_0000000000000001;               // addi $8, $6, 1 (loop2)
            memory[45] <= 32'b001000_10001_01010_0000000000000000;               // lw $10, 0($17)
            memory[46] <= 32'b010101_00000000000000000000000000;                 // syscall
            memory[47] <= 32'b000001_10010_10010_0000000000000001;               // addi $18, $18, 1
            memory[48] <= 32'b000001_10001_10001_0000000000000001;               // addi $17, $17, 1
            memory[49] <= 32'b001011_11011_10010_1111111111111010;               // bne $18, $27, -6
            memory[50] <= 32'b010001_00000000000000000000010000;                 // jr $16 (end2)
            cur <= 51;
        end
    end
    
    // Sequential write operation at posedge of clk.
    always @(posedge reset or posedge clk) begin
        if(reset==1'b1) begin
            dataout <= 0;
            for(i=cur;i<depth;i=i+1) begin memory[i] <= 0; end
        end
        else begin
            if(writeEnable==1'b1 && mode==1'b0) begin
                memory[address_a] <= in;
            end
        end
    end

    // Combinational read operation.
    assign out = memory[address_b];
endmodule


/// This is the module which will be used as the source of memory and this has the following controls as explained
// clk - The synchronizing signal for all the phases of the processor machine.
// reset - The reset signal to delete and restart the whole memory.
// in - The data which is send as input for storing in memory.
// out - The data which is being asked for from memory.
// mode - The working mode of the memory currently. 0 means write mode and 1 means read only mode.
// address_a - The address at which the input is filled by the memory.
// address_b - The address from which output is generated by the memory.
// writeEnable - In write mode when we have to refrain from writing into memory disable this flag.
module veda_data #(parameter width = 32, parameter depth = 256, parameter len = 8, parameter start = 0) (
    clk,reset,
    in,out,mode,address_a,address_b,
    writeEnable
);
    input wire [width-1:0] in;
    input wire [len-1:0] address_a,address_b;
    input wire clk,reset,mode,writeEnable;                            // Mode 0 means write mode and Mode 1 means read mode
    output wire [width-1:0] out;
    
    reg [width-1:0] memory[0:depth-1];
    reg [width-1:0] dataout,cur;
    integer i;

    // Setting the memory at erased state.
    initial begin
        if(start == 0) begin cur <= 0; end
    end
    
    // Load the default data of bubble sort if start is set to HIGH.
    initial begin
        if(start == 1) begin
            // Write program to enter data memory into the machine
            memory[0]  <= " ";                           // strCT
            memory[1]  <= "\n";                          // strCR
            memory[2]  <= "Init";                        // strInit
            memory[3]  <= "ial ";
            memory[4]  <= "arra";
            memory[5]  <= "y:  ";
            memory[6]  <= "Sort";                        // strResult
            memory[7]  <= "ed a";
            memory[8]  <= "rray";
            memory[9]  <= ":   ";
            memory[10] <= 32'd11;                        // n
            memory[11] <= 32'd643;                       // arr
            memory[12] <= 32'd573;
            memory[13] <= 32'd532;
            memory[14] <= 32'd087;
            memory[15] <= 32'd879;
            memory[16] <= 32'd242;
            memory[17] <= 32'd64;
            memory[18] <= 32'd805;
            memory[19] <= 32'd868;
            memory[20] <= 32'd57320;
            memory[21] <= 32'd378;
            cur <= 22;
        end
    end
    
    // Sequential write operation at posedge of clk.
    always @(posedge reset or posedge clk) begin
        if(reset==1'b1) begin
            dataout <= 0;
            for(i=cur;i<depth;i=i+1) begin memory[i] <= 0; end
        end
        else begin
            if(writeEnable==1'b1 && mode==1'b0) begin
                memory[address_a] <= in;
            end
        end
    end

    // Combinational read operation.
    assign out = memory[address_b];
endmodule
